library ieee;
use ieee.std_logic_1164.all;


package reg_file_port is

    constant REG_R0 : std_logic_vector(2 downto 0) := "000";
    constant REG_R1 : std_logic_vector(2 downto 0) := "001";
    constant REG_R2 : std_logic_vector(2 downto 0) := "010";
    constant REG_R3 : std_logic_vector(2 downto 0) := "011";
    constant REG_R4 : std_logic_vector(2 downto 0) := "100";
    constant REG_R5 : std_logic_vector(2 downto 0) := "101";
    constant REG_R6 : std_logic_vector(2 downto 0) := "110";
    constant REG_R7 : std_logic_vector(2 downto 0) := "111";

end package reg_file_port;


---------------------------------------------------------------------------------
-- MIT License
--
-- Copyright (c) 2015-2018 Dominik Salvet
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.
---------------------------------------------------------------------------------
