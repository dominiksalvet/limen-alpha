library ieee;
use ieee.std_logic_1164.all;


package limen_alpha_public is
    
    constant CORE_0_INT_ADDR   : std_ulogic_vector(15 downto 0) := x"0004";
    constant CORE_0_IP_REG_RST : std_ulogic_vector(15 downto 0) := x"0000";
    constant CORE_0_PRNG_SEED  : std_ulogic_vector(15 downto 0) := x"ffff";
    
    constant CORE_1_INT_ADDR   : std_ulogic_vector(15 downto 0) := x"000c";
    constant CORE_1_IP_REG_RST : std_ulogic_vector(15 downto 0) := x"0008";
    constant CORE_1_PRNG_SEED  : std_ulogic_vector(15 downto 0) := x"ddd4";
    
end package limen_alpha_public;


--------------------------------------------------------------------------------
-- MIT License
--
-- Copyright (c) 2018 Dominik Salvet
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.
--------------------------------------------------------------------------------
